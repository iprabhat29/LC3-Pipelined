module mon(lc3Interface.MONITOR inf);

endmodule